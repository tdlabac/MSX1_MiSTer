module msx1
(
	input         clk,
	input         reset
);

endmodule
